module gray_count(
                input           clk,
                input           enable,
                input           reset_L,
                input   [4:0]   count,
                output  [4:0]   salida_gray );




endmodule
